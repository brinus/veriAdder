module ADDER ( input    [24:0] WORD_0,
                        [24:0] WORD_1,
                        [24:0] WORD_2,
                        [24:0] WORD_3,
                        [24:0] WORD_4,
                        [24:0] WORD_5,
                        [24:0] WORD_6,
                        [24:0] WORD_7,
                        [24:0] WORD_8,
                        [24:0] WORD_9,
                        [24:0] WORD_10,
                        [24:0] WORD_11,
                        [24:0] WORD_12,
                        [24:0] WORD_13,
                        [24:0] WORD_14,
                        [24:0] WORD_15,
                        CLK,
                output  [24:0] RES);

                always @ (posedge CLK) begin
                               
                end
endmodule