`ifndef _global_parameters_vh
`define _global_parameters_vh

`define LYCALOQBIT      25
`define NSERDESBP       16
`define LYBOARDS        16

`endif