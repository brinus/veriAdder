module ADDER_TB ();

endmodule